`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 		David Brown
//// 
//// Create Date:    12/3/2025 
//// Module Name:    vgaGlyphRom
//// Project Name: 	vga
//// Description: 	
////
//// Dependencies: 	
////
//// Revision 0.01 - File Created
////
////////////////////////////////////////////////////////////////////////////////////
//
//
//////////////////////////////////////////////////////////////////////////////////

module vgaGlyphRom(clk,  address, q);

input clk;
input [13:0]address;

output reg [7:0] q;

reg [7:0] rom [0:16383];

initial begin
    $readmemh("font8x8.hex", rom);
end

always @(posedge clk)
    q <= rom[address];

endmodule